** Generated for: hspiceD
** Generated on: Apr 22 22:52:21 2015
** Design library name: ECE8893_lib
** Design cell name: abat_invchain_latched
** Design view name: schematic
.PARAM c=0.2525m


.TRAN 10e-9 5e-6 START=0.0
.OPTION DELMAX=10e-9


.OP

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/nethome/jshinsato3/ECE6130_Cadence/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_nom/PMOS_VTL.inc"
.INCLUDE "/nethome/jshinsato3/ECE6130_Cadence/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_nom/PMOS_VTH.inc"
.INCLUDE "/nethome/jshinsato3/ECE6130_Cadence/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_nom/PMOS_VTG.inc"
.INCLUDE "/nethome/jshinsato3/ECE6130_Cadence/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_nom/PMOS_THKOX.inc"
.INCLUDE "/nethome/jshinsato3/ECE6130_Cadence/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_nom/NMOS_VTL.inc"
.INCLUDE "/nethome/jshinsato3/ECE6130_Cadence/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_nom/NMOS_VTH.inc"
.INCLUDE "/nethome/jshinsato3/ECE6130_Cadence/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_nom/NMOS_VTG.inc"
.INCLUDE "/nethome/jshinsato3/ECE6130_Cadence/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_nom/NMOS_THKOX.inc"

** Library name: ECE8893_lib
** Cell name: nand2
** View name: schematic
.subckt nand2 a b out vground vsupply
m1 out a vsupply vsupply PMOS_VTH L=45e-9 W=360e-9
m0 out b vsupply vsupply PMOS_VTH L=45e-9 W=360e-9
m3 net22 b vground vground NMOS_VTH L=45e-9 W=157.5e-9
m2 out a net22 vground NMOS_VTH L=45e-9 W=157.5e-9
.ends nand2
** End of subcircuit definition.

** Library name: ECE8893_lib
** Cell name: inv1
** View name: schematic
.subckt inv1 a out vground vsupply
m1 out a vsupply vsupply PMOS_VTH L=45e-9 W=360e-9
m3 out a vground vground NMOS_VTH L=45e-9 W=90e-9
.ends inv1
** End of subcircuit definition.

** Library name: ECE8893_lib
** Cell name: abat_latch
** View name: schematic
.subckt abat_latch clk d q q__ vsupply vground
xi3 net12 q__ q vground vsupply nand2
xi2 q net15 q__ vground vsupply nand2
xi1 clk net17 net15 vground vsupply nand2
xi0 d clk net12 vground vsupply nand2
xi5 d net17 vground vsupply inv1
.ends abat_latch
** End of subcircuit definition.

** Library name: ECE8893_lib
** Cell name: abat_invchain_latched
** View name: schematic
r1 vcc net130 1e-9
r0 v1 net131 1e-9
xi1 vcc chain_out q q__ vccdc vss abat_latch
c1 net130 vss 'c*1e-3'
c0 net131 vss 'c*1e-3'
l1 vref vcc 1e-6
l0 v1 vref 1e-6
m22 vcc v1 vss vss NMOS_VTG L=45e-9 W=90e-9
m20 vss vcc v1 vss NMOS_VTG L=45e-9 W=180e-9
m23 vcc v1 vccdc vccdc PMOS_VTG L=45e-9 W=90e-9
m21 vccdc vcc v1 vccdc PMOS_VTG L=45e-9 W=180e-9
m18 chain_out net121 vss 0 NMOS_VTH L=45e-9 W=1.77147e-3
m16 net121 net118 vss 0 NMOS_VTH L=45e-9 W=590.49e-6
m15 net118 net114 vss 0 NMOS_VTH L=45e-9 W=196.83e-6
m12 net114 net110 vss 0 NMOS_VTH L=45e-9 W=65.61e-6
m10 net110 net107 vss 0 NMOS_VTH L=45e-9 W=21.87e-6
m8 net107 net104 vss 0 NMOS_VTH L=45e-9 W=7.29e-6
m7 net104 net101 vss 0 NMOS_VTH L=45e-9 W=2.43e-6
m4 net101 net96 vss 0 NMOS_VTH L=45e-9 W=810e-9
m2 net96 net89 vss 0 NMOS_VTH L=45e-9 W=270e-9
m0 net89 in vss 0 NMOS_VTH L=45e-9 W=90e-9
m19 chain_out net121 vcc vcc PMOS_VTH L=45e-9 W=2.36196e-3
m17 net121 net118 vcc vcc PMOS_VTH L=45e-9 W=787.32e-6
m14 net118 net114 vcc vcc PMOS_VTH L=45e-9 W=262.44e-6
m13 net114 net110 vcc vcc PMOS_VTH L=45e-9 W=87.48e-6
m11 net110 net107 vcc vcc PMOS_VTH L=45e-9 W=29.16e-6
m9 net107 net104 vcc vcc PMOS_VTH L=45e-9 W=9.72e-6
m6 net104 net101 vcc vcc PMOS_VTH L=45e-9 W=3.24e-6
m5 net101 net96 vcc vcc PMOS_VTH L=45e-9 W=1.08e-6
m3 net96 net89 vcc vcc PMOS_VTH L=45e-9 W=360e-9
m1 net89 in vcc vcc PMOS_VTH L=45e-9 W=360e-9
.include "/nethome/jshinsato3/simulation/abat_invchain_latched/hspiceD/schematic/netlist/_graphical_stimuli.scs"
.END
